
library IEEE; 
use IEEE.STD_LOGIC_1164.all; 
use STD.TEXTIO.all;
use IEEE.NUMERIC_STD.all; 

entity dmem is -- data memory
  port(clk, we:  in STD_LOGIC;
       a, wd:    in STD_LOGIC_VECTOR(31 downto 0);
       rd:       out STD_LOGIC_VECTOR(31 downto 0));
end;

architecture behave of dmem is
	type ramtype is array (63 downto 0) of STD_LOGIC_VECTOR(31 downto 0);
	signal mem: ramtype;
begin
	process(clk)
	begin
		if clk'event and clk = '1' then
			if we = '1' then	mem(to_integer(unsigned(a))) <= wd;
			end if;
			
			rd <= mem(to_integer(unsigned(a)));
		end if;
	end process;
end;
